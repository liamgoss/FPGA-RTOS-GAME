// GameSystem.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module GameSystem (
		input  wire        clk_clk,            //         clk.clk
		input  wire [2:0]  keys_export,        //        keys.export
		inout  wire [7:0]  lcd_DATA,           //         lcd.DATA
		output wire        lcd_ON,             //            .ON
		output wire        lcd_BLON,           //            .BLON
		output wire        lcd_EN,             //            .EN
		output wire        lcd_RS,             //            .RS
		output wire        lcd_RW,             //            .RW
		output wire [7:0]  ledg_export,        //        ledg.export
		output wire [17:0] leds_export,        //        leds.export
		input  wire        reset_reset_n,      //       reset.reset_n
		output wire [12:0] sdram_wire_addr,    //  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,      //            .ba
		output wire        sdram_wire_cas_n,   //            .cas_n
		output wire        sdram_wire_cke,     //            .cke
		output wire        sdram_wire_cs_n,    //            .cs_n
		inout  wire [31:0] sdram_wire_dq,      //            .dq
		output wire [3:0]  sdram_wire_dqm,     //            .dqm
		output wire        sdram_wire_ras_n,   //            .ras_n
		output wire        sdram_wire_we_n,    //            .we_n
		output wire [6:0]  seven_seg_0_export, // seven_seg_0.export
		output wire [6:0]  seven_seg_1_export, // seven_seg_1.export
		output wire [6:0]  seven_seg_2_export, // seven_seg_2.export
		output wire [6:0]  seven_seg_3_export, // seven_seg_3.export
		output wire [6:0]  seven_seg_4_export, // seven_seg_4.export
		output wire [6:0]  seven_seg_5_export, // seven_seg_5.export
		output wire [6:0]  seven_seg_6_export, // seven_seg_6.export
		output wire [6:0]  seven_seg_7_export, // seven_seg_7.export
		input  wire [17:0] switches_export     //    switches.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_lcd_avalon_lcd_slave_chipselect;           // mm_interconnect_0:lcd_avalon_lcd_slave_chipselect -> lcd:chipselect
	wire   [7:0] mm_interconnect_0_lcd_avalon_lcd_slave_readdata;             // lcd:readdata -> mm_interconnect_0:lcd_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest;          // lcd:waitrequest -> mm_interconnect_0:lcd_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_lcd_avalon_lcd_slave_address;              // mm_interconnect_0:lcd_avalon_lcd_slave_address -> lcd:address
	wire         mm_interconnect_0_lcd_avalon_lcd_slave_read;                 // mm_interconnect_0:lcd_avalon_lcd_slave_read -> lcd:read
	wire         mm_interconnect_0_lcd_avalon_lcd_slave_write;                // mm_interconnect_0:lcd_avalon_lcd_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_0_lcd_avalon_lcd_slave_writedata;            // mm_interconnect_0:lcd_avalon_lcd_slave_writedata -> lcd:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                      // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                       // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_ledg_s1_chipselect;                        // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                          // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                           // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_write;                             // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                         // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_keys_s1_chipselect;                        // mm_interconnect_0:KEYS_s1_chipselect -> KEYS:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                          // KEYS:readdata -> mm_interconnect_0:KEYS_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                           // mm_interconnect_0:KEYS_s1_address -> KEYS:address
	wire         mm_interconnect_0_keys_s1_write;                             // mm_interconnect_0:KEYS_s1_write -> KEYS:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                         // mm_interconnect_0:KEYS_s1_writedata -> KEYS:writedata
	wire         mm_interconnect_0_seven_seg_0_s1_chipselect;                 // mm_interconnect_0:seven_seg_0_s1_chipselect -> seven_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_readdata;                   // seven_seg_0:readdata -> mm_interconnect_0:seven_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_0_s1_address;                    // mm_interconnect_0:seven_seg_0_s1_address -> seven_seg_0:address
	wire         mm_interconnect_0_seven_seg_0_s1_write;                      // mm_interconnect_0:seven_seg_0_s1_write -> seven_seg_0:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_writedata;                  // mm_interconnect_0:seven_seg_0_s1_writedata -> seven_seg_0:writedata
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                 // mm_interconnect_0:seven_seg_1_s1_chipselect -> seven_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                   // seven_seg_1:readdata -> mm_interconnect_0:seven_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                    // mm_interconnect_0:seven_seg_1_s1_address -> seven_seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                      // mm_interconnect_0:seven_seg_1_s1_write -> seven_seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                  // mm_interconnect_0:seven_seg_1_s1_writedata -> seven_seg_1:writedata
	wire         mm_interconnect_0_seven_seg_2_s1_chipselect;                 // mm_interconnect_0:seven_seg_2_s1_chipselect -> seven_seg_2:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_readdata;                   // seven_seg_2:readdata -> mm_interconnect_0:seven_seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_2_s1_address;                    // mm_interconnect_0:seven_seg_2_s1_address -> seven_seg_2:address
	wire         mm_interconnect_0_seven_seg_2_s1_write;                      // mm_interconnect_0:seven_seg_2_s1_write -> seven_seg_2:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_writedata;                  // mm_interconnect_0:seven_seg_2_s1_writedata -> seven_seg_2:writedata
	wire         mm_interconnect_0_seven_seg_3_s1_chipselect;                 // mm_interconnect_0:seven_seg_3_s1_chipselect -> seven_seg_3:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_readdata;                   // seven_seg_3:readdata -> mm_interconnect_0:seven_seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_3_s1_address;                    // mm_interconnect_0:seven_seg_3_s1_address -> seven_seg_3:address
	wire         mm_interconnect_0_seven_seg_3_s1_write;                      // mm_interconnect_0:seven_seg_3_s1_write -> seven_seg_3:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_writedata;                  // mm_interconnect_0:seven_seg_3_s1_writedata -> seven_seg_3:writedata
	wire         mm_interconnect_0_seven_seg_5_s1_chipselect;                 // mm_interconnect_0:seven_seg_5_s1_chipselect -> seven_seg_5:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_readdata;                   // seven_seg_5:readdata -> mm_interconnect_0:seven_seg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_5_s1_address;                    // mm_interconnect_0:seven_seg_5_s1_address -> seven_seg_5:address
	wire         mm_interconnect_0_seven_seg_5_s1_write;                      // mm_interconnect_0:seven_seg_5_s1_write -> seven_seg_5:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_writedata;                  // mm_interconnect_0:seven_seg_5_s1_writedata -> seven_seg_5:writedata
	wire         mm_interconnect_0_seven_seg_4_s1_chipselect;                 // mm_interconnect_0:seven_seg_4_s1_chipselect -> seven_seg_4:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_readdata;                   // seven_seg_4:readdata -> mm_interconnect_0:seven_seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_4_s1_address;                    // mm_interconnect_0:seven_seg_4_s1_address -> seven_seg_4:address
	wire         mm_interconnect_0_seven_seg_4_s1_write;                      // mm_interconnect_0:seven_seg_4_s1_write -> seven_seg_4:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_writedata;                  // mm_interconnect_0:seven_seg_4_s1_writedata -> seven_seg_4:writedata
	wire         mm_interconnect_0_seven_seg_6_s1_chipselect;                 // mm_interconnect_0:seven_seg_6_s1_chipselect -> seven_seg_6:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_6_s1_readdata;                   // seven_seg_6:readdata -> mm_interconnect_0:seven_seg_6_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_6_s1_address;                    // mm_interconnect_0:seven_seg_6_s1_address -> seven_seg_6:address
	wire         mm_interconnect_0_seven_seg_6_s1_write;                      // mm_interconnect_0:seven_seg_6_s1_write -> seven_seg_6:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_6_s1_writedata;                  // mm_interconnect_0:seven_seg_6_s1_writedata -> seven_seg_6:writedata
	wire         mm_interconnect_0_system_timer_s1_chipselect;                // mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                  // system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                   // mm_interconnect_0:system_timer_s1_address -> system_timer:address
	wire         mm_interconnect_0_system_timer_s1_write;                     // mm_interconnect_0:system_timer_s1_write -> system_timer:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                 // mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;              // mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                // high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                 // mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_0_high_res_timer_s1_write;                   // mm_interconnect_0:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;               // mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_seven_seg_7_s1_chipselect;                 // mm_interconnect_0:seven_seg_7_s1_chipselect -> seven_seg_7:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_7_s1_readdata;                   // seven_seg_7:readdata -> mm_interconnect_0:seven_seg_7_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_7_s1_address;                    // mm_interconnect_0:seven_seg_7_s1_address -> seven_seg_7:address
	wire         mm_interconnect_0_seven_seg_7_s1_write;                      // mm_interconnect_0:seven_seg_7_s1_write -> seven_seg_7:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_7_s1_writedata;                  // mm_interconnect_0:seven_seg_7_s1_writedata -> seven_seg_7:writedata
	wire         irq_mapper_receiver0_irq;                                    // KEYS:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // system_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // high_res_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [KEYS:reset_n, high_res_timer:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, lcd:reset, ledg:reset_n, leds:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sdram:reset_n, seven_seg_0:reset_n, seven_seg_1:reset_n, seven_seg_2:reset_n, seven_seg_3:reset_n, seven_seg_4:reset_n, seven_seg_5:reset_n, seven_seg_6:reset_n, seven_seg_7:reset_n, switches:reset_n, sysid_qsys_0:reset_n, system_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> onchip_memory2_0:reset_req

	GameSystem_KEYS keys (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_export),                          // external_connection.export
		.irq        (irq_mapper_receiver0_irq)              //                 irq.irq
	);

	GameSystem_high_res_timer high_res_timer (
		.clk        (clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                        //   irq.irq
	);

	GameSystem_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                     //               irq.irq
	);

	GameSystem_lcd lcd (
		.clk         (clk_clk),                                            //                clk.clk
		.reset       (rst_controller_reset_out_reset),                     //              reset.reset
		.address     (mm_interconnect_0_lcd_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_lcd_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_lcd_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_lcd_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_lcd_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_lcd_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_DATA),                                           // external_interface.export
		.LCD_ON      (lcd_ON),                                             //                   .export
		.LCD_BLON    (lcd_BLON),                                           //                   .export
		.LCD_EN      (lcd_EN),                                             //                   .export
		.LCD_RS      (lcd_RS),                                             //                   .export
		.LCD_RW      (lcd_RW)                                              //                   .export
	);

	GameSystem_ledg ledg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	GameSystem_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	GameSystem_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	GameSystem_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	GameSystem_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	GameSystem_seven_seg_0 seven_seg_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_0_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_0_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_2_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_2_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_3_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_3_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_4_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_4_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_5_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_5_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_6_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_6_export)                           // external_connection.export
	);

	GameSystem_seven_seg_0 seven_seg_7 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_7_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_7_export)                           // external_connection.export
	);

	GameSystem_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	GameSystem_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	GameSystem_system_timer system_timer (
		.clk        (clk_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                      //   irq.irq
	);

	GameSystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                     //                                     clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                              //      nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                    (nios2_gen2_0_data_master_address),                            //                      nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                (nios2_gen2_0_data_master_waitrequest),                        //                                              .waitrequest
		.nios2_gen2_0_data_master_byteenable                 (nios2_gen2_0_data_master_byteenable),                         //                                              .byteenable
		.nios2_gen2_0_data_master_read                       (nios2_gen2_0_data_master_read),                               //                                              .read
		.nios2_gen2_0_data_master_readdata                   (nios2_gen2_0_data_master_readdata),                           //                                              .readdata
		.nios2_gen2_0_data_master_readdatavalid              (nios2_gen2_0_data_master_readdatavalid),                      //                                              .readdatavalid
		.nios2_gen2_0_data_master_write                      (nios2_gen2_0_data_master_write),                              //                                              .write
		.nios2_gen2_0_data_master_writedata                  (nios2_gen2_0_data_master_writedata),                          //                                              .writedata
		.nios2_gen2_0_data_master_debugaccess                (nios2_gen2_0_data_master_debugaccess),                        //                                              .debugaccess
		.nios2_gen2_0_instruction_master_address             (nios2_gen2_0_instruction_master_address),                     //               nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest         (nios2_gen2_0_instruction_master_waitrequest),                 //                                              .waitrequest
		.nios2_gen2_0_instruction_master_read                (nios2_gen2_0_instruction_master_read),                        //                                              .read
		.nios2_gen2_0_instruction_master_readdata            (nios2_gen2_0_instruction_master_readdata),                    //                                              .readdata
		.nios2_gen2_0_instruction_master_readdatavalid       (nios2_gen2_0_instruction_master_readdatavalid),               //                                              .readdatavalid
		.high_res_timer_s1_address                           (mm_interconnect_0_high_res_timer_s1_address),                 //                             high_res_timer_s1.address
		.high_res_timer_s1_write                             (mm_interconnect_0_high_res_timer_s1_write),                   //                                              .write
		.high_res_timer_s1_readdata                          (mm_interconnect_0_high_res_timer_s1_readdata),                //                                              .readdata
		.high_res_timer_s1_writedata                         (mm_interconnect_0_high_res_timer_s1_writedata),               //                                              .writedata
		.high_res_timer_s1_chipselect                        (mm_interconnect_0_high_res_timer_s1_chipselect),              //                                              .chipselect
		.jtag_uart_0_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                 jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                              .write
		.jtag_uart_0_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                              .read
		.jtag_uart_0_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                              .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                              .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                              .chipselect
		.KEYS_s1_address                                     (mm_interconnect_0_keys_s1_address),                           //                                       KEYS_s1.address
		.KEYS_s1_write                                       (mm_interconnect_0_keys_s1_write),                             //                                              .write
		.KEYS_s1_readdata                                    (mm_interconnect_0_keys_s1_readdata),                          //                                              .readdata
		.KEYS_s1_writedata                                   (mm_interconnect_0_keys_s1_writedata),                         //                                              .writedata
		.KEYS_s1_chipselect                                  (mm_interconnect_0_keys_s1_chipselect),                        //                                              .chipselect
		.lcd_avalon_lcd_slave_address                        (mm_interconnect_0_lcd_avalon_lcd_slave_address),              //                          lcd_avalon_lcd_slave.address
		.lcd_avalon_lcd_slave_write                          (mm_interconnect_0_lcd_avalon_lcd_slave_write),                //                                              .write
		.lcd_avalon_lcd_slave_read                           (mm_interconnect_0_lcd_avalon_lcd_slave_read),                 //                                              .read
		.lcd_avalon_lcd_slave_readdata                       (mm_interconnect_0_lcd_avalon_lcd_slave_readdata),             //                                              .readdata
		.lcd_avalon_lcd_slave_writedata                      (mm_interconnect_0_lcd_avalon_lcd_slave_writedata),            //                                              .writedata
		.lcd_avalon_lcd_slave_waitrequest                    (mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest),          //                                              .waitrequest
		.lcd_avalon_lcd_slave_chipselect                     (mm_interconnect_0_lcd_avalon_lcd_slave_chipselect),           //                                              .chipselect
		.ledg_s1_address                                     (mm_interconnect_0_ledg_s1_address),                           //                                       ledg_s1.address
		.ledg_s1_write                                       (mm_interconnect_0_ledg_s1_write),                             //                                              .write
		.ledg_s1_readdata                                    (mm_interconnect_0_ledg_s1_readdata),                          //                                              .readdata
		.ledg_s1_writedata                                   (mm_interconnect_0_ledg_s1_writedata),                         //                                              .writedata
		.ledg_s1_chipselect                                  (mm_interconnect_0_ledg_s1_chipselect),                        //                                              .chipselect
		.leds_s1_address                                     (mm_interconnect_0_leds_s1_address),                           //                                       leds_s1.address
		.leds_s1_write                                       (mm_interconnect_0_leds_s1_write),                             //                                              .write
		.leds_s1_readdata                                    (mm_interconnect_0_leds_s1_readdata),                          //                                              .readdata
		.leds_s1_writedata                                   (mm_interconnect_0_leds_s1_writedata),                         //                                              .writedata
		.leds_s1_chipselect                                  (mm_interconnect_0_leds_s1_chipselect),                        //                                              .chipselect
		.nios2_gen2_0_debug_mem_slave_address                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                  nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                              .write
		.nios2_gen2_0_debug_mem_slave_read                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                              .read
		.nios2_gen2_0_debug_mem_slave_readdata               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                              .readdata
		.nios2_gen2_0_debug_mem_slave_writedata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                              .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                              .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                              .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                              .debugaccess
		.onchip_memory2_0_s1_address                         (mm_interconnect_0_onchip_memory2_0_s1_address),               //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                           (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                              .write
		.onchip_memory2_0_s1_readdata                        (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                              .readdata
		.onchip_memory2_0_s1_writedata                       (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                              .writedata
		.onchip_memory2_0_s1_byteenable                      (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                              .byteenable
		.onchip_memory2_0_s1_chipselect                      (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                              .chipselect
		.onchip_memory2_0_s1_clken                           (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                              .clken
		.sdram_s1_address                                    (mm_interconnect_0_sdram_s1_address),                          //                                      sdram_s1.address
		.sdram_s1_write                                      (mm_interconnect_0_sdram_s1_write),                            //                                              .write
		.sdram_s1_read                                       (mm_interconnect_0_sdram_s1_read),                             //                                              .read
		.sdram_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                         //                                              .readdata
		.sdram_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                        //                                              .writedata
		.sdram_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                       //                                              .byteenable
		.sdram_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                              .readdatavalid
		.sdram_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                      //                                              .waitrequest
		.sdram_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect),                       //                                              .chipselect
		.seven_seg_0_s1_address                              (mm_interconnect_0_seven_seg_0_s1_address),                    //                                seven_seg_0_s1.address
		.seven_seg_0_s1_write                                (mm_interconnect_0_seven_seg_0_s1_write),                      //                                              .write
		.seven_seg_0_s1_readdata                             (mm_interconnect_0_seven_seg_0_s1_readdata),                   //                                              .readdata
		.seven_seg_0_s1_writedata                            (mm_interconnect_0_seven_seg_0_s1_writedata),                  //                                              .writedata
		.seven_seg_0_s1_chipselect                           (mm_interconnect_0_seven_seg_0_s1_chipselect),                 //                                              .chipselect
		.seven_seg_1_s1_address                              (mm_interconnect_0_seven_seg_1_s1_address),                    //                                seven_seg_1_s1.address
		.seven_seg_1_s1_write                                (mm_interconnect_0_seven_seg_1_s1_write),                      //                                              .write
		.seven_seg_1_s1_readdata                             (mm_interconnect_0_seven_seg_1_s1_readdata),                   //                                              .readdata
		.seven_seg_1_s1_writedata                            (mm_interconnect_0_seven_seg_1_s1_writedata),                  //                                              .writedata
		.seven_seg_1_s1_chipselect                           (mm_interconnect_0_seven_seg_1_s1_chipselect),                 //                                              .chipselect
		.seven_seg_2_s1_address                              (mm_interconnect_0_seven_seg_2_s1_address),                    //                                seven_seg_2_s1.address
		.seven_seg_2_s1_write                                (mm_interconnect_0_seven_seg_2_s1_write),                      //                                              .write
		.seven_seg_2_s1_readdata                             (mm_interconnect_0_seven_seg_2_s1_readdata),                   //                                              .readdata
		.seven_seg_2_s1_writedata                            (mm_interconnect_0_seven_seg_2_s1_writedata),                  //                                              .writedata
		.seven_seg_2_s1_chipselect                           (mm_interconnect_0_seven_seg_2_s1_chipselect),                 //                                              .chipselect
		.seven_seg_3_s1_address                              (mm_interconnect_0_seven_seg_3_s1_address),                    //                                seven_seg_3_s1.address
		.seven_seg_3_s1_write                                (mm_interconnect_0_seven_seg_3_s1_write),                      //                                              .write
		.seven_seg_3_s1_readdata                             (mm_interconnect_0_seven_seg_3_s1_readdata),                   //                                              .readdata
		.seven_seg_3_s1_writedata                            (mm_interconnect_0_seven_seg_3_s1_writedata),                  //                                              .writedata
		.seven_seg_3_s1_chipselect                           (mm_interconnect_0_seven_seg_3_s1_chipselect),                 //                                              .chipselect
		.seven_seg_4_s1_address                              (mm_interconnect_0_seven_seg_4_s1_address),                    //                                seven_seg_4_s1.address
		.seven_seg_4_s1_write                                (mm_interconnect_0_seven_seg_4_s1_write),                      //                                              .write
		.seven_seg_4_s1_readdata                             (mm_interconnect_0_seven_seg_4_s1_readdata),                   //                                              .readdata
		.seven_seg_4_s1_writedata                            (mm_interconnect_0_seven_seg_4_s1_writedata),                  //                                              .writedata
		.seven_seg_4_s1_chipselect                           (mm_interconnect_0_seven_seg_4_s1_chipselect),                 //                                              .chipselect
		.seven_seg_5_s1_address                              (mm_interconnect_0_seven_seg_5_s1_address),                    //                                seven_seg_5_s1.address
		.seven_seg_5_s1_write                                (mm_interconnect_0_seven_seg_5_s1_write),                      //                                              .write
		.seven_seg_5_s1_readdata                             (mm_interconnect_0_seven_seg_5_s1_readdata),                   //                                              .readdata
		.seven_seg_5_s1_writedata                            (mm_interconnect_0_seven_seg_5_s1_writedata),                  //                                              .writedata
		.seven_seg_5_s1_chipselect                           (mm_interconnect_0_seven_seg_5_s1_chipselect),                 //                                              .chipselect
		.seven_seg_6_s1_address                              (mm_interconnect_0_seven_seg_6_s1_address),                    //                                seven_seg_6_s1.address
		.seven_seg_6_s1_write                                (mm_interconnect_0_seven_seg_6_s1_write),                      //                                              .write
		.seven_seg_6_s1_readdata                             (mm_interconnect_0_seven_seg_6_s1_readdata),                   //                                              .readdata
		.seven_seg_6_s1_writedata                            (mm_interconnect_0_seven_seg_6_s1_writedata),                  //                                              .writedata
		.seven_seg_6_s1_chipselect                           (mm_interconnect_0_seven_seg_6_s1_chipselect),                 //                                              .chipselect
		.seven_seg_7_s1_address                              (mm_interconnect_0_seven_seg_7_s1_address),                    //                                seven_seg_7_s1.address
		.seven_seg_7_s1_write                                (mm_interconnect_0_seven_seg_7_s1_write),                      //                                              .write
		.seven_seg_7_s1_readdata                             (mm_interconnect_0_seven_seg_7_s1_readdata),                   //                                              .readdata
		.seven_seg_7_s1_writedata                            (mm_interconnect_0_seven_seg_7_s1_writedata),                  //                                              .writedata
		.seven_seg_7_s1_chipselect                           (mm_interconnect_0_seven_seg_7_s1_chipselect),                 //                                              .chipselect
		.switches_s1_address                                 (mm_interconnect_0_switches_s1_address),                       //                                   switches_s1.address
		.switches_s1_readdata                                (mm_interconnect_0_switches_s1_readdata),                      //                                              .readdata
		.sysid_qsys_0_control_slave_address                  (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //                    sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                 (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                              .readdata
		.system_timer_s1_address                             (mm_interconnect_0_system_timer_s1_address),                   //                               system_timer_s1.address
		.system_timer_s1_write                               (mm_interconnect_0_system_timer_s1_write),                     //                                              .write
		.system_timer_s1_readdata                            (mm_interconnect_0_system_timer_s1_readdata),                  //                                              .readdata
		.system_timer_s1_writedata                           (mm_interconnect_0_system_timer_s1_writedata),                 //                                              .writedata
		.system_timer_s1_chipselect                          (mm_interconnect_0_system_timer_s1_chipselect)                 //                                              .chipselect
	);

	GameSystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
